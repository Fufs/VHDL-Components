LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY  IS
  port(  : IN ; 
     : OUT );
END ;

ARCHITECTURE struct OF  IS
BEGIN
  
END struct;